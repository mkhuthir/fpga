// Muthanna Alwahash
// (c) Sept 2023

module ()


endmodule